`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:19:56 03/02/2025
// Design Name:   Pipeline
// Module Name:   E:/Documents and Settings/student/EE533_Lab7/EE533_Lab_7/Pipeline_tb.v
// Project Name:  EE533_Lab_7
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Pipeline
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Pipeline_tb;

	// Inputs
	reg clk;
	reg [31:0] Instr_IN;
	reg Instr_W_en;
	reg [8:0] I_W_Addr;
	reg [63:0] ONE;
	reg rst;

	// Outputs
	wire ADDI_EX;
	wire ADDI_ID;
	wire ADDI_M;
	wire ADDI_WB;
	wire [63:0] ALU_B;
	wire [3:0] ALU_OP_EX;
	wire [3:0] ALU_OP_ID;
	wire [63:0] ALU_result_EX;
	wire [63:0] ALU_result_M;
	wire [63:0] ALU_result_WB;
	wire BEQ_ID;
	wire BGT_ID;
	wire BLT_ID;
	wire [7:0] D_MEM_addr;
	wire [63:0] D_out_M;
	wire [63:0] D_out_WB;
	wire [31:0] Instruction;
	wire J_ID;
	wire LW_EX;
	wire LW_ID;
	wire LW_M;
	wire LW_WB;
	wire MOVI_EX;
	wire MOVI_ID;
	wire MOVI_M;
	wire MOVI_WB;
	wire NOOP_EX;
	wire NOOP_ID;
	wire NOOP_M;
	wire NOOP_WB;
	wire [63:0] Offset_EX;
	wire [63:0] Offset_ID;
	wire [63:0] Offset_M;
	wire [63:0] Offset_WB;
	wire [5:0] OP_CODE_ID;
	wire [63:0] PC;
	wire PC_ctrl;
	wire [63:0] PC_next;
	wire [63:0] PC_plus_one;
	wire [63:0] RF_WB_Din;
	wire [63:0] rs_data_EX;
	wire [63:0] rs_data_ID;
	wire [63:0] rs_data_M;
	wire [63:0] rs_data_WB;
	wire [4:0] rs_ID;
	wire [63:0] rt_data_EX;
	wire [63:0] rt_data_ID;
	wire [63:0] rt_data_M;
	wire [4:0] rt_EX;
	wire [4:0] rt_ID;
	wire [4:0] rt_M;
	wire [2:0] rt_WB;
	wire SW_EX;
	wire SW_ID;
	wire SW_M;
	wire SW_WB;
	wire WME_EX;
	wire WME_ID;
	wire WME_M;
	wire WRE_EX;
	wire WRE_ID;
	wire WRE_M;
	wire WRE_WB;

	// Instantiate the Unit Under Test (UUT)
	Pipeline uut (
		.clk(clk), 
		.Instr_IN(Instr_IN), 
		.Instr_W_en(Instr_W_en), 
		.I_W_Addr(I_W_Addr), 
		.ONE(ONE), 
		.rst(rst), 
		.ADDI_EX(ADDI_EX), 
		.ADDI_ID(ADDI_ID), 
		.ADDI_M(ADDI_M), 
		.ADDI_WB(ADDI_WB), 
		.ALU_B(ALU_B), 
		.ALU_OP_EX(ALU_OP_EX), 
		.ALU_OP_ID(ALU_OP_ID), 
		.ALU_result_EX(ALU_result_EX), 
		.ALU_result_M(ALU_result_M), 
		.ALU_result_WB(ALU_result_WB), 
		.BEQ_ID(BEQ_ID), 
		.BGT_ID(BGT_ID), 
		.BLT_ID(BLT_ID), 
		.D_MEM_addr(D_MEM_addr), 
		.D_out_M(D_out_M), 
		.D_out_WB(D_out_WB), 
		.Instruction(Instruction), 
		.J_ID(J_ID), 
		.LW_EX(LW_EX), 
		.LW_ID(LW_ID), 
		.LW_M(LW_M), 
		.LW_WB(LW_WB), 
		.MOVI_EX(MOVI_EX), 
		.MOVI_ID(MOVI_ID), 
		.MOVI_M(MOVI_M), 
		.MOVI_WB(MOVI_WB), 
		.NOOP_EX(NOOP_EX), 
		.NOOP_ID(NOOP_ID), 
		.NOOP_M(NOOP_M), 
		.NOOP_WB(NOOP_WB), 
		.Offset_EX(Offset_EX), 
		.Offset_ID(Offset_ID), 
		.Offset_M(Offset_M), 
		.Offset_WB(Offset_WB), 
		.OP_CODE_ID(OP_CODE_ID), 
		.PC(PC), 
		.PC_ctrl(PC_ctrl), 
		.PC_next(PC_next), 
		.PC_plus_one(PC_plus_one), 
		.RF_WB_Din(RF_WB_Din), 
		.rs_data_EX(rs_data_EX), 
		.rs_data_ID(rs_data_ID), 
		.rs_data_M(rs_data_M), 
		.rs_data_WB(rs_data_WB), 
		.rs_ID(rs_ID), 
		.rt_data_EX(rt_data_EX), 
		.rt_data_ID(rt_data_ID), 
		.rt_data_M(rt_data_M), 
		.rt_EX(rt_EX), 
		.rt_ID(rt_ID), 
		.rt_M(rt_M), 
		.rt_WB(rt_WB), 
		.SW_EX(SW_EX), 
		.SW_ID(SW_ID), 
		.SW_M(SW_M), 
		.SW_WB(SW_WB), 
		.WME_EX(WME_EX), 
		.WME_ID(WME_ID), 
		.WME_M(WME_M), 
		.WRE_EX(WRE_EX), 
		.WRE_ID(WRE_ID), 
		.WRE_M(WRE_M), 
		.WRE_WB(WRE_WB)
	);

	always #50 clk = ~clk;

	initial begin
		// Initialize Inputs
		clk = 1;
		Instr_IN = 0;
		Instr_W_en = 0;
		I_W_Addr = 0;
		ONE = 0;
		rst = 1;

		// Wait 100 ns for global reset to finish
		@(posedge clk);
		ONE = 64'd1;
		rst = 0;
        
		// Add stimulus here
		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);

		@(posedge clk);
		$stop;

	end
      
endmodule

